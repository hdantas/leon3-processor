library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_arith.all; 
use ieee.std_logic_unsigned.all;

entity qSelector is
	port (
		signed	: in std_logic;
		x     	: in  std_logic_vector(64 downto 0);
		d     	: in  std_logic_vector(31 downto 0);
		q    	: out std_logic_vector(2 downto 0)
	);
end;

architecture rtl of qSelector is

type qgen_lut_t is array ( 0 to 255) of std_logic_vector(2 downto 0);
--Index => d[k-1..k-5] & x[2k-1..2k-5]
constant qgen_lut: qgen_lut_t := (
	136 => "011",		--10001000
	137 => "011",		--10001001
	138 => "011",		--10001010
	139 => "010",		--10001011
	140 => "010",		--10001100
	141 => "001",		--10001101
	142 => "001",		--10001110
	143 => "000",		--10001111
	128 => "000",		--10000000
	129 => "111",		--10000001
	130 => "111",		--10000010
	131 => "110",		--10000011
	132 => "110",		--10000100
	133 => "101",		--10000101
	134 => "101",		--10000110
	135 => "101",		--10000111
	152 => "---",		--10011000
	153 => "011",		--10011001
	154 => "011",		--10011010
	155 => "011",		--10011011
	156 => "010",		--10011100
	157 => "001",		--10011101
	158 => "001",		--10011110
	159 => "000",		--10011111
	144 => "000",		--10010000
	145 => "111",		--10010001
	146 => "111",		--10010010
	147 => "110",		--10010011
	148 => "101",		--10010100
	149 => "101",		--10010101
	150 => "101",		--10010110
	151 => "---",		--10010111
	168 => "---",		--10101000
	169 => "---",		--10101001
	170 => "011",		--10101010
	171 => "011",		--10101011
	172 => "011",		--10101100
	173 => "010",		--10101101
	174 => "001",		--10101110
	175 => "000",		--10101111
	160 => "000",		--10100000
	161 => "111",		--10100001
	162 => "110",		--10100010
	163 => "101",		--10100011
	164 => "101",		--10100100
	165 => "101",		--10100101
	166 => "---",		--10100110
	167 => "---",		--10100111
	184 => "---",		--10111000
	185 => "---",		--10111001
	186 => "---",		--10111010
	187 => "011",		--10111011
	188 => "011",		--10111100
	189 => "010",		--10111101
	190 => "001",		--10111110
	191 => "000",		--10111111
	176 => "000",		--10110000
	177 => "111",		--10110001
	178 => "110",		--10110010
	179 => "101",		--10110011
	180 => "101",		--10110100
	181 => "---",		--10110101
	182 => "---",		--10110110
	183 => "---",		--10110111
	200 => "---",		--11001000
	201 => "---",		--11001001
	202 => "---",		--11001010
	203 => "---",		--11001011
	204 => "---",		--11001100
	205 => "---",		--11001101
	206 => "---",		--11001110
	207 => "---",		--11001111
	192 => "---",		--11000000
	193 => "---",		--11000001
	194 => "---",		--11000010
	195 => "---",		--11000011
	196 => "---",		--11000100
	197 => "---",		--11000101
	198 => "---",		--11000110
	199 => "---",		--11000111
	216 => "---",		--11011000
	217 => "---",		--11011001
	218 => "---",		--11011010
	219 => "---",		--11011011
	220 => "---",		--11011100
	221 => "---",		--11011101
	222 => "---",		--11011110
	223 => "---",		--11011111
	208 => "---",		--11010000
	209 => "---",		--11010001
	210 => "---",		--11010010
	211 => "---",		--11010011
	212 => "---",		--11010100
	213 => "---",		--11010101
	214 => "---",		--11010110
	215 => "---",		--11010111
	232 => "---",		--11101000
	233 => "---",		--11101001
	234 => "---",		--11101010
	235 => "---",		--11101011
	236 => "---",		--11101100
	237 => "---",		--11101101
	238 => "---",		--11101110
	239 => "---",		--11101111
	224 => "---",		--11100000
	225 => "---",		--11100001
	226 => "---",		--11100010
	227 => "---",		--11100011
	228 => "---",		--11100100
	229 => "---",		--11100101
	230 => "---",		--11100110
	231 => "---",		--11100111
	248 => "---",		--11111000
	249 => "---",		--11111001
	250 => "---",		--11111010
	251 => "---",		--11111011
	252 => "---",		--11111100
	253 => "---",		--11111101
	254 => "---",		--11111110
	255 => "---",		--11111111
	240 => "---",		--11110000
	241 => "---",		--11110001
	242 => "---",		--11110010
	243 => "---",		--11110011
	244 => "---",		--11110100
	245 => "---",		--11110101
	246 => "---",		--11110110
	247 => "---",		--11110111
	8 => "---",		--00001000
	9 => "---",		--00001001
	10 => "---",		--00001010
	11 => "---",		--00001011
	12 => "---",		--00001100
	13 => "---",		--00001101
	14 => "---",		--00001110
	15 => "---",		--00001111
	0 => "---",		--00000000
	1 => "---",		--00000001
	2 => "---",		--00000010
	3 => "---",		--00000011
	4 => "---",		--00000100
	5 => "---",		--00000101
	6 => "---",		--00000110
	7 => "---",		--00000111
	24 => "---",		--00011000
	25 => "---",		--00011001
	26 => "---",		--00011010
	27 => "---",		--00011011
	28 => "---",		--00011100
	29 => "---",		--00011101
	30 => "---",		--00011110
	31 => "---",		--00011111
	16 => "---",		--00010000
	17 => "---",		--00010001
	18 => "---",		--00010010
	19 => "---",		--00010011
	20 => "---",		--00010100
	21 => "---",		--00010101
	22 => "---",		--00010110
	23 => "---",		--00010111
	40 => "---",		--00101000
	41 => "---",		--00101001
	42 => "---",		--00101010
	43 => "---",		--00101011
	44 => "---",		--00101100
	45 => "---",		--00101101
	46 => "---",		--00101110
	47 => "---",		--00101111
	32 => "---",		--00100000
	33 => "---",		--00100001
	34 => "---",		--00100010
	35 => "---",		--00100011
	36 => "---",		--00100100
	37 => "---",		--00100101
	38 => "---",		--00100110
	39 => "---",		--00100111
	56 => "---",		--00111000
	57 => "---",		--00111001
	58 => "---",		--00111010
	59 => "---",		--00111011
	60 => "---",		--00111100
	61 => "---",		--00111101
	62 => "---",		--00111110
	63 => "---",		--00111111
	48 => "---",		--00110000
	49 => "---",		--00110001
	50 => "---",		--00110010
	51 => "---",		--00110011
	52 => "---",		--00110100
	53 => "---",		--00110101
	54 => "---",		--00110110
	55 => "---",		--00110111
	72 => "---",		--01001000
	73 => "---",		--01001001
	74 => "---",		--01001010
	75 => "101",		--01001011
	76 => "101",		--01001100
	77 => "110",		--01001101
	78 => "111",		--01001110
	79 => "111",		--01001111
	64 => "000",		--01000000
	65 => "001",		--01000001
	66 => "010",		--01000010
	67 => "011",		--01000011
	68 => "011",		--01000100
	69 => "---",		--01000101
	70 => "---",		--01000110
	71 => "---",		--01000111
	88 => "---",		--01011000
	89 => "---",		--01011001
	90 => "101",		--01011010
	91 => "101",		--01011011
	92 => "101",		--01011100
	93 => "110",		--01011101
	94 => "111",		--01011110
	95 => "000",		--01011111
	80 => "000",		--01010000
	81 => "001",		--01010001
	82 => "010",		--01010010
	83 => "011",		--01010011
	84 => "011",		--01010100
	85 => "011",		--01010101
	86 => "---",		--01010110
	87 => "---",		--01010111
	104 => "---",		--01101000
	105 => "101",		--01101001
	106 => "101",		--01101010
	107 => "101",		--01101011
	108 => "110",		--01101100
	109 => "110",		--01101101
	110 => "111",		--01101110
	111 => "000",		--01101111
	96 => "000",		--01100000
	97 => "001",		--01100001
	98 => "001",		--01100010
	99 => "010",		--01100011
	100 => "011",		--01100100
	101 => "011",		--01100101
	102 => "011",		--01100110
	103 => "---",		--01100111
	120 => "101",		--01111000
	121 => "101",		--01111001
	122 => "101",		--01111010
	123 => "110",		--01111011
	124 => "110",		--01111100
	125 => "111",		--01111101
	126 => "111",		--01111110
	127 => "000",		--01111111
	112 => "000",		--01110000
	113 => "001",		--01110001
	114 => "001",		--01110010
	115 => "010",		--01110011
	116 => "010",		--01110100
	117 => "011",		--01110101
	118 => "011",		--01110110
	119 => "011"		--01110111
);

begin
  process(x(63 downto 0),d)
    begin
		if (x="1110000000000000000000000000000000000000000000000000000000000000") and (d="01000000000000000000000000000000") then
			q<="110";
		elsif (x="1101000000000000000000000000000000000000000000000000000000000000") and (d="01000000000000000000000000000000") then
			q<="101";
		else
			if(signed='1') then
				q<=qgen_lut(conv_integer(d(31 downto 28) & x(63 downto 60)));
				--q<="000";
			else
				q<=qgen_lut(conv_integer('0' & d(31 downto 29) & x(64 downto 61)));
			end if;
		end if;		
	end process;
end;