library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_arith.all; 
use ieee.std_logic_unsigned.all;

entity qSelector is
	port (
		signed	: in std_logic;
		x     	: in  std_logic_vector(64 downto 0);
		d     	: in  std_logic_vector(31 downto 0);
		q    	: out std_logic_vector(2 downto 0)
	);
end;

architecture rtl of qSelector is

type qgen_lut_t is array ( 0 to 127) of std_logic_vector(2 downto 0);
--Index => d[k-2..k-5] & x[2k-1..2k-5]
constant qgen_lut : qgen_lut_t := (
	8 => "---",			--0001000
	9 => "---",			--0001001
	10 => "---",		--0001010
	11 => "---",		--0001011
	12 => "---",		--0001100
	13 => "---",		--0001101
	14 => "---",		--0001110
	15 => "---",		--0001111
	0 => "---",			--0000000
	1 => "---",			--0000001
	2 => "---",			--0000010
	3 => "---",			--0000011
	4 => "---",			--0000100
	5 => "---",			--0000101
	6 => "---",			--0000110
	7 => "---",			--0000111
	24 => "---",		--0011000
	25 => "---",		--0011001
	26 => "---",		--0011010
	27 => "---",		--0011011
	28 => "---",		--0011100
	29 => "---",		--0011101
	30 => "---",		--0011110
	31 => "---",		--0011111
	16 => "---",		--0010000
	17 => "---",		--0010001
	18 => "---",		--0010010
	19 => "---",		--0010011
	20 => "---",		--0010100
	21 => "---",		--0010101
	22 => "---",		--0010110
	23 => "---",		--0010111
	40 => "---",		--0101000
	41 => "---",		--0101001
	42 => "---",		--0101010
	43 => "---",		--0101011
	44 => "---",		--0101100
	45 => "---",		--0101101
	46 => "---",		--0101110
	47 => "---",		--0101111
	32 => "---",		--0100000
	33 => "---",		--0100001
	34 => "---",		--0100010
	35 => "---",		--0100011
	36 => "---",		--0100100
	37 => "---",		--0100101
	38 => "---",		--0100110
	39 => "---",		--0100111
	56 => "---",		--0111000
	57 => "---",		--0111001
	58 => "---",		--0111010
	59 => "---",		--0111011
	60 => "---",		--0111100
	61 => "---",		--0111101
	62 => "---",		--0111110
	63 => "---",		--0111111
	48 => "---",		--0110000
	49 => "---",		--0110001
	50 => "---",		--0110010
	51 => "---",		--0110011
	52 => "---",		--0110100
	53 => "---",		--0110101
	54 => "---",		--0110110
	55 => "---",		--0110111
	72 => "---",		--1001000
	73 => "---",		--1001001
	74 => "---",		--1001010
	75 => "101",		--1001011
	76 => "101",		--1001100
	77 => "110",		--1001101
	78 => "111",		--1001110
	79 => "111",		--1001111
	64 => "000",		--1000000
	65 => "001",		--1000001
	66 => "010",		--1000010
	67 => "011",		--1000011
	68 => "011",		--1000100
	69 => "---",		--1000101
	70 => "---",		--1000110
	71 => "---",		--1000111
	88 => "---",		--1011000
	89 => "---",		--1011001
	90 => "101",		--1011010
	91 => "101",		--1011011
	92 => "101",		--1011100
	93 => "110",		--1011101
	94 => "111",		--1011110
	95 => "000",		--1011111
	80 => "000",		--1010000
	81 => "001",		--1010001
	82 => "010",		--1010010
	83 => "011",		--1010011
	84 => "011",		--1010100
	85 => "011",		--1010101
	86 => "---",		--1010110
	87 => "---",		--1010111
	104 => "---",		--1101000
	105 => "101",		--1101001
	106 => "101",		--1101010
	107 => "101",		--1101011
	108 => "110",		--1101100
	109 => "110",		--1101101
	110 => "111",		--1101110
	111 => "000",		--1101111
	96 => "000",		--1100000
	97 => "001",		--1100001
	98 => "001",		--1100010
	99 => "010",		--1100011
	100 => "011",		--1100100
	101 => "011",		--1100101
	102 => "011",		--1100110
	103 => "---",		--1100111
	120 => "101",		--1111000
	121 => "101",		--1111001
	122 => "101",		--1111010
	123 => "110",		--1111011
	124 => "110",		--1111100
	125 => "111",		--1111101
	126 => "111",		--1111110
	127 => "000",		--1111111
	112 => "000",		--1110000
	113 => "001",		--1110001
	114 => "001",		--1110010
	115 => "010",		--1110011
	116 => "010",		--1110100
	117 => "011",		--1110101
	118 => "011",		--1110110
	119 => "011"		--1110111
);

begin
  process(x(63 downto 0),d)
    begin
		if (x="1110000000000000000000000000000000000000000000000000000000000000") and (d="01000000000000000000000000000000") then
			q<="110";
		elsif (x="1101000000000000000000000000000000000000000000000000000000000000") and (d="01000000000000000000000000000000") then
			q<="101";
		else
			if(signed='1') then
				q<=qgen_lut(conv_integer(d(30 downto 28) & x(63 downto 60)));
				--q<="000";
			else
				q<=qgen_lut(conv_integer(d(31 downto 29) & x(64 downto 61)));
			end if;
		end if;		
	end process;
end;