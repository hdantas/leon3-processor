/home/nuno/repos/pdp/Multiplier/src/mul32_3cycle.vhd