#
# Automatically generated make config: don't edit
#

#
# Synthesis      
#
# CONFIG_SYN_INFERRED is not set
# CONFIG_SYN_STRATIX is not set
# CONFIG_SYN_STRATIXII is not set
# CONFIG_SYN_STRATIXIII is not set
# CONFIG_SYN_CYCLONEIII is not set
# CONFIG_SYN_ALTERA is not set
# CONFIG_SYN_AXCEL is not set
# CONFIG_SYN_PROASIC is not set
# CONFIG_SYN_PROASICPLUS is not set
# CONFIG_SYN_PROASIC3 is not set
# CONFIG_SYN_UT025CRH is not set
# CONFIG_SYN_ATC18 is not set
# CONFIG_SYN_ATC18RHA is not set
# CONFIG_SYN_CUSTOM1 is not set
# CONFIG_SYN_EASIC90 is not set
# CONFIG_SYN_IHP25 is not set
# CONFIG_SYN_IHP25RH is not set
# CONFIG_SYN_LATTICE is not set
# CONFIG_SYN_ECLIPSE is not set
# CONFIG_SYN_PEREGRINE is not set
# CONFIG_SYN_RH_LIB18T is not set
# CONFIG_SYN_RHUMC is not set
# CONFIG_SYN_SMIC13 is not set
# CONFIG_SYN_SPARTAN2 is not set
# CONFIG_SYN_SPARTAN3 is not set
# CONFIG_SYN_SPARTAN3E is not set
# CONFIG_SYN_VIRTEX is not set
# CONFIG_SYN_VIRTEXE is not set
# CONFIG_SYN_VIRTEX2 is not set
CONFIG_SYN_VIRTEX4=y
# CONFIG_SYN_VIRTEX5 is not set
# CONFIG_SYN_UMC is not set
# CONFIG_SYN_TSMC90 is not set
# CONFIG_SYN_INFER_RAM is not set
# CONFIG_SYN_INFER_PADS is not set
# CONFIG_SYN_NO_ASYNC is not set
# CONFIG_SYN_SCAN is not set

#
# Clock generation
#
# CONFIG_CLK_INFERRED is not set
# CONFIG_CLK_HCLKBUF is not set
# CONFIG_CLK_ALTDLL is not set
# CONFIG_CLK_LATDLL is not set
# CONFIG_CLK_PRO3PLL is not set
# CONFIG_CLK_LIB18T is not set
# CONFIG_CLK_RHUMC is not set
# CONFIG_CLK_CLKDLL is not set
CONFIG_CLK_DCM=y
CONFIG_CLK_MUL=16
CONFIG_CLK_DIV=20
# CONFIG_PCI_CLKDLL is not set
# CONFIG_CLK_NOFB is not set
# CONFIG_PCI_SYSCLK is not set
CONFIG_LEON3=y
CONFIG_PROC_NUM=1

#
# Processor            
#

#
# Integer unit                                           
#
CONFIG_IU_NWINDOWS=8
CONFIG_IU_V8MULDIV=y
# CONFIG_IU_MUL_LATENCY_2 is not set
# CONFIG_IU_MUL_LATENCY_4 is not set
CONFIG_IU_MUL_LATENCY_5=y
# CONFIG_IU_MUL_MAC is not set
CONFIG_IU_SVT=y
CONFIG_IU_LDELAY=1
CONFIG_IU_WATCHPOINTS=1
CONFIG_PWD=y
CONFIG_IU_RSTADDR=00000

#
# Floating-point unit
#
# CONFIG_FPU_ENABLE is not set

#
# Cache system
#
CONFIG_ICACHE_ENABLE=y
# CONFIG_ICACHE_ASSO1 is not set
CONFIG_ICACHE_ASSO2=y
# CONFIG_ICACHE_ASSO3 is not set
# CONFIG_ICACHE_ASSO4 is not set
# CONFIG_ICACHE_SZ1 is not set
# CONFIG_ICACHE_SZ2 is not set
# CONFIG_ICACHE_SZ4 is not set
CONFIG_ICACHE_SZ8=y
# CONFIG_ICACHE_SZ16 is not set
# CONFIG_ICACHE_SZ32 is not set
# CONFIG_ICACHE_SZ64 is not set
# CONFIG_ICACHE_SZ128 is not set
# CONFIG_ICACHE_SZ256 is not set
# CONFIG_ICACHE_LZ16 is not set
CONFIG_ICACHE_LZ32=y
# CONFIG_ICACHE_ALGORND is not set
CONFIG_ICACHE_ALGOLRR=y
# CONFIG_ICACHE_ALGOLRU is not set
# CONFIG_ICACHE_LOCK is not set
CONFIG_DCACHE_ENABLE=y
# CONFIG_DCACHE_ASSO1 is not set
CONFIG_DCACHE_ASSO2=y
# CONFIG_DCACHE_ASSO3 is not set
# CONFIG_DCACHE_ASSO4 is not set
# CONFIG_DCACHE_SZ1 is not set
# CONFIG_DCACHE_SZ2 is not set
CONFIG_DCACHE_SZ4=y
# CONFIG_DCACHE_SZ8 is not set
# CONFIG_DCACHE_SZ16 is not set
# CONFIG_DCACHE_SZ32 is not set
# CONFIG_DCACHE_SZ64 is not set
# CONFIG_DCACHE_SZ128 is not set
# CONFIG_DCACHE_SZ256 is not set
CONFIG_DCACHE_LZ16=y
# CONFIG_DCACHE_LZ32 is not set
# CONFIG_DCACHE_ALGORND is not set
CONFIG_DCACHE_ALGOLRR=y
# CONFIG_DCACHE_ALGOLRU is not set
# CONFIG_DCACHE_LOCK is not set
CONFIG_DCACHE_SNOOP=y
# CONFIG_DCACHE_SNOOP_FAST is not set
# CONFIG_DCACHE_SNOOP_SEPTAG is not set
CONFIG_CACHE_FIXED=0

#
# MMU
#
CONFIG_MMU_ENABLE=y
CONFIG_MMU_COMBINED=y
# CONFIG_MMU_SPLIT is not set
# CONFIG_MMU_REPARRAY is not set
CONFIG_MMU_REPINCREMENT=y
# CONFIG_MMU_I2 is not set
# CONFIG_MMU_I4 is not set
CONFIG_MMU_I8=y
# CONFIG_MMU_I16 is not set
# CONFIG_MMU_I32 is not set

#
# Debug Support Unit        
#
CONFIG_DSU_ENABLE=y
CONFIG_DSU_ITRACE=y
# CONFIG_DSU_ITRACESZ1 is not set
CONFIG_DSU_ITRACESZ2=y
# CONFIG_DSU_ITRACESZ4 is not set
# CONFIG_DSU_ITRACESZ8 is not set
# CONFIG_DSU_ITRACESZ16 is not set
CONFIG_DSU_ATRACE=y
# CONFIG_DSU_ATRACESZ1 is not set
CONFIG_DSU_ATRACESZ2=y
# CONFIG_DSU_ATRACESZ4 is not set
# CONFIG_DSU_ATRACESZ8 is not set
# CONFIG_DSU_ATRACESZ16 is not set

#
# Fault-tolerance  
#

#
# VHDL debug settings       
#
# CONFIG_IU_DISAS is not set
# CONFIG_DEBUG_PC32 is not set

#
# AMBA configuration
#
CONFIG_AHB_DEFMST=0
CONFIG_AHB_RROBIN=y
# CONFIG_AHB_SPLIT is not set
CONFIG_AHB_IOADDR=FFF
CONFIG_APB_HADDR=800
# CONFIG_AHB_MON is not set

#
# Debug Link           
#
CONFIG_DSU_UART=y
CONFIG_DSU_JTAG=y

#
# Peripherals             
#

#
# Memory controller             
#

#
# Leon2 memory controller        
#
CONFIG_MCTRL_LEON2=y
# CONFIG_MCTRL_8BIT is not set
# CONFIG_MCTRL_16BIT is not set
# CONFIG_MCTRL_5CS is not set
# CONFIG_MCTRL_SDRAM is not set

#
# DDR266 SDRAM controller             
#
CONFIG_DDRSP=y
CONFIG_DDRSP_INIT=y
CONFIG_DDRSP_FREQ=100
CONFIG_DDRSP_COL=9
CONFIG_DDRSP_MBYTE=64
CONFIG_DDRSP_RSKEW=0

#
# Synchronous SRAM controller   
#
# CONFIG_SSCTRL is not set
CONFIG_AHBSTAT_ENABLE=y
CONFIG_AHBSTAT_NFTSLV=1

#
# On-chip RAM/ROM                 
#
# CONFIG_AHBROM_ENABLE is not set
# CONFIG_AHBRAM_ENABLE is not set

#
# Ethernet             
#
# CONFIG_GRETH_ENABLE is not set

#
# UART, timer, I2C, I/O port and interrupt controller
#
CONFIG_UART1_ENABLE=y
# CONFIG_UA1_FIFO1 is not set
# CONFIG_UA1_FIFO2 is not set
CONFIG_UA1_FIFO4=y
# CONFIG_UA1_FIFO8 is not set
# CONFIG_UA1_FIFO16 is not set
# CONFIG_UA1_FIFO32 is not set
CONFIG_IRQ3_ENABLE=y
# CONFIG_IRQ3_SEC is not set
CONFIG_GPT_ENABLE=y
CONFIG_GPT_NTIM=2
CONFIG_GPT_SW=8
CONFIG_GPT_TW=32
CONFIG_GPT_IRQ=8
CONFIG_GPT_SEPIRQ=y
# CONFIG_GPT_WDOGEN is not set
CONFIG_GRGPIO_ENABLE=y
CONFIG_GRGPIO_WIDTH=14
CONFIG_GRGPIO_IMASK=0FFFE
# CONFIG_I2C_ENABLE is not set

#
# Keybord and VGA interface
#
# CONFIG_KBD_ENABLE is not set
# CONFIG_VGA_ENABLE is not set
# CONFIG_SVGA_ENABLE is not set

#
# VHDL Debugging        
#
# CONFIG_DEBUG_UART is not set
