/home/nuno/repos/pdp/Multiplier/src/mul32_1cycle.vhd